interface dut_if(input logic clk);
  logic       rst_n;
  logic [7:0] a;
  logic [7:0] b;
  logic [8:0] y;
endinterface
