package tb_pkg;
  `include "uvm_macros.svh"
  `include "uvm_transaction.sv"
  `include "uvm_driver.sv"
  `include "uvm_monitor.sv"
  `include "uvm_scoreboard.sv"
  `include "uvm_env.sv"
  `include "uvm_sequence.sv"
  `include "uvm_test.sv"
  import uvm_pkg::*;

endpackage